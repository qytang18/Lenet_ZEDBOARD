`ifndef _define_header_vh_
`define _define_header_vh_

// state_index
`define IDLE  0
`define SCONV_1  1
`define SPOOL_1 2
`define SCONV_2 3
`define SPOOL_2 4
`define SFC_1 5
`define SFC_2 6
`define SFC_3 7

// parameter
`define MAC_NUM 120
`define MAX_NUM 15
`endif