`ifndef _define_header_vh_
`define _define_header_vh_

// state_index
`define IDLE  0
`define SCONV_1  1
`define SPOOL_1 2
`define SCONV_2 3
`define SPOOL_2 4
`define SFC_1 5
`define SRELU_1 6
`define SFC_2 7
`define SRELU_2 8
`define SFC_3 9

// parameter
`define MAC_NUM 120
`define MAX_NUM 15
`endif